module async_rom_case
    ( 
      input  wire  [7:0] r_addr,
      output reg  [28:0] r_data
    );


    // body
    always @*
        case (r_addr)
				// Fetch
            8'h00 : r_data = 29'b00000000100001000000010110101;
            8'h01 : r_data = 29'b00000000000001000000010000000;
            8'h02 : r_data = 29'b01100000000010000000010000000;
            8'h03 : r_data = 29'b00000000000000100000010000000;
            8'h04 : r_data = 29'b00000000000000010001011000000;//sin interrupcion
				
            8'h05 : r_data = 29'b00000000000000101000010000000;
            8'h06 : r_data = 29'b01100000100110000010010000000;
            8'h07 : r_data = 29'b00010010000010000001111000000;
				
				//mov ACC, A
            8'h08 : r_data = 29'b10000001111110000001111000000;
            8'h09 : r_data = 29'b00000000000000000000000000000;//desde aqui no se usan
            8'h0A : r_data = 29'b00000000000000000000000000000;
            8'h0B : r_data = 29'b00000000000000000000000000000;
            8'h0C : r_data = 29'b00000000000000000000000000000;
            8'h0D : r_data = 29'b00000000000000000000000000000;
            8'h0E : r_data = 29'b00000000000000000000000000000;
            8'h0F : r_data = 29'b00000000000000000000000000000;
				
				//mov A, ACCC                   //Intclr
            8'h10 : r_data = 29'b10000011101110000001111000000;
            8'h11 : r_data = 29'b00000000000000000000000000000;
            8'h12 : r_data = 29'b00000000000000000000000000000;
            8'h13 : r_data = 29'b00000000000000000000000000000;
            8'h14 : r_data = 29'b00000000000000000000000000000;
            8'h15 : r_data = 29'b00000000000000000000000000000;
            8'h16 : r_data = 29'b00000000000000000000000000000;
            8'h17 : r_data = 29'b00000000000000000000000000000;
				
				
				
				//mov ACC, CTE
				
				8'h18 : r_data = 29'b00000000000001000000010000000;
            8'h19 : r_data = 29'b01100000000010000000010000000;
            8'h1A : r_data = 29'b00000000000000110000010000000;
            8'h1B : r_data = 29'b00000000011110010001111000000;
            8'h1C : r_data = 29'b00000000000000000000000000000;
            8'h1D : r_data = 29'b00000000000000000000000000000;
            8'h1E : r_data = 29'b00000000000000000000000000000;
            8'h1F : r_data = 29'b00000000000000000000000000000;
				
				
				//mov ACC,[DPTR]   ---YA ESTA EN LAS DIAPOS
            8'h20 : r_data = 29'b00000001000001000000010000000;
            8'h21 : r_data = 29'b00000000000000000000010000000;
            8'h22 : r_data = 29'b00000000000000100000010000000;
            8'h23 : r_data = 29'b00000000011110010001111000000;
            8'h24 : r_data = 29'b00000000000000000000000000000;
            8'h25 : r_data = 29'b00000000000000000000000000000;
            8'h26 : r_data = 29'b00000000000000000000000000000;
            8'h27 : r_data = 29'b00000000000000000000000000000;
				
				//MOV DPTR, ACC   --REVISAR          ------------------
				
            8'h28 : r_data = 29'b10000011101010000001111000000;
            8'h29 : r_data = 29'b00000000000000000000000000000;
            8'h2A : r_data = 29'b00000000000000000000000000000;
            8'h2B : r_data = 29'b00000000000000000000000000000;
            8'h2C : r_data = 29'b00000000000000000000000000000;
            8'h2D : r_data = 29'b00000000000000000000000000000;
            8'h2E : r_data = 29'b00000000000000000000000000000;
            8'h2F : r_data = 29'b00000000000000000000000000000;
				
				
				//MOC [DPTR],ACC   --REVISAR                ------------
            8'h30 : r_data = 29'b10000001000001000000010000000;
            8'h31 : r_data = 29'b10000011100000100000010000000;
            8'h32 : r_data = 29'b10000000001000000011111000000;
            8'h33 : r_data = 29'b00000000000000000000000000000;
            8'h34 : r_data = 29'b00000000000000000000000000000;
            8'h35 : r_data = 29'b00000000000000000000000000000;
            8'h36 : r_data = 29'b00000000000000000000000000000;
            8'h37 : r_data = 29'b00000000000000000000000000000;
				
				//INV ACC
            8'h38 : r_data = 29'b10010011111110100001111000000;
            8'h39 : r_data = 29'b00000000000000000000000000000;
            8'h3A : r_data = 29'b00000000000000000000000000000;
            8'h3B : r_data = 29'b00000000000000000000000000000;
            8'h3C : r_data = 29'b00000000000000000000000000000;
            8'h3D : r_data = 29'b00000000000000000000000000000;
            8'h3E : r_data = 29'b00000000000000000000000000000;
            8'h3F : r_data = 29'b00000000000000000000000000000;
				
				//AND ACC, A
				
            8'h40 : r_data = 29'b10100001111110100001111000000;
            8'h41 : r_data = 29'b00000000000000000000000000000;
            8'h42 : r_data = 29'b00000000000000000000000000000;
            8'h43 : r_data = 29'b00000000000000000000000000000;
            8'h44 : r_data = 29'b00000000000000000000000000000;
            8'h45 : r_data = 29'b00000000000000000000000000000;
            8'h46 : r_data = 29'b00000000000000000000000000000;
            8'h47 : r_data = 29'b00000000000000000000000000000;
				
				//ADD ACC, A   //revisar nuestro vs profe
					
            8'h48 : r_data = 29'b11010001111110000000101000000;
            8'h49 : r_data = 29'b00000000000000000000000000000;
            8'h4A : r_data = 29'b00000000000000000000000000000;
            8'h4B : r_data = 29'b00000000000000000000000000000;
            8'h4C : r_data = 29'b00000000000000000000000000000;
            8'h4D : r_data = 29'b00000000000000000000000000000;
            8'h4E : r_data = 29'b00000000000000000000000000000;
            8'h4F : r_data = 29'b00000000000000000000000000000;
				
				//JMP DIR  --REVISARRRRRRRRRRR              ------------
				
            8'h50 : r_data = 29'b00000000000001000000010001010;
            8'h51 : r_data = 29'b01100000000010000001111000000;
            8'h52 : r_data = 29'b00000000000000000000010000000;
            8'h53 : r_data = 29'b00000000000000100000010000000;
            8'h54 : r_data = 29'b00000000000010010001111000000;
            8'h55 : r_data = 29'b00000000000010010001111000000;
            8'h56 : r_data = 29'b00000000000000000000000000000;
            8'h57 : r_data = 29'b00000000000000000000000000000;
				
				//JZ DIR   --REVISAR                        -------------
				
            8'h58 : r_data = 29'b00000000000001000000010010010;
            8'h59 : r_data = 29'b01100000000010000001111000000;
            8'h5A : r_data = 29'b00000000000000000000010000000;
            8'h5B : r_data = 29'b00000000000000100000010000000;
            8'h5C : r_data = 29'b00000000000010010001111000000;
            8'h5D : r_data = 29'b00000000000010010001111000000;
            8'h5E : r_data = 29'b00000000000000000000000000000;
            8'h5F : r_data = 29'b00000000000000000000000000000;
            
				
				//JN DIR  

				8'h60 : r_data = 29'b00000000000001000000010011010;
            8'h61 : r_data = 29'b01100000000010000001111000000;
            8'h62 : r_data = 29'b00000000000000000000010000000;
            8'h63 : r_data = 29'b00000000000000100000010000000;
            8'h64 : r_data = 29'b00000000000010010001111000000;
            8'h65 : r_data = 29'b00000000000010010001111000000;
            8'h66 : r_data = 29'b00000000000000000000000000000;
            8'h67 : r_data = 29'b00000000000000000000000000000;
				
				//JC DIR
				
				8'h68 : r_data = 29'b00000000000001000000010100010;
            8'h69 : r_data = 29'b01100000000010000001111000000;
            8'h6A : r_data = 29'b00000000000000000000010000000;
            8'h6B : r_data = 29'b00000000000000100000010000000;
            8'h6C : r_data = 29'b00000000000010010001111000000;
            8'h6D : r_data = 29'b00000000000010010001111000000;
            8'h6E : r_data = 29'b00000000000000000000000000000;
            8'h6F : r_data = 29'b00000000000000000000000000000;
				
				//CALL DIR                   --revisarrrr --------------  
            8'h70 : r_data = 29'b00000000000000000000000000000;
            8'h71 : r_data = 29'b00000000000000000000000000000;
            8'h72 : r_data = 29'b00000000000000000000000000000;
            8'h73 : r_data = 29'b00000000000000000000000000000;
            8'h74 : r_data = 29'b00000000000000000000000000000;
            8'h75 : r_data = 29'b00000000000000000000000000000;
            8'h76 : r_data = 29'b00000000000000000000000000000;
            8'h77 : r_data = 29'b00000000000000000000000000000;
				
				//RET                           ---revisar preguntarrrr
            8'h78 : r_data = 29'b00000000000000000000000000000; 
            8'h79 : r_data = 29'b00000000000000000000000000000;
            8'h7A : r_data = 29'b00000000000000000000000000000;
            8'h7B : r_data = 29'b00000000000000000000000000000;
            8'h7C : r_data = 29'b00000000000000000000000000000;
            8'h7D : r_data = 29'b00000000000000000000000000000;
            8'h7E : r_data = 29'b00000000000000000000000000000;
            8'h7F : r_data = 29'b00000000000000000000000000000;
				
				//OR ACC, A ---------------------------------------------------------------retomar desde aqui
            8'h80 : r_data = 29'b10110001111110100001111000000;
            8'h81 : r_data = 29'b00000000000000000000000000000;
            8'h82 : r_data = 29'b00000000000000000000000000000;
            8'h83 : r_data = 29'b00000000000000000000000000000;
            8'h84 : r_data = 29'b00000000000000000000000000000;
            8'h85 : r_data = 29'b00000000000000000000000000000;
            8'h86 : r_data = 29'b00000000000000000000000000000;
            8'h87 : r_data = 29'b00000000000000000000000000000;
				
				//XOR ACC,A
            8'h88 : r_data = 29'b11000001111110100001111000000;
            8'h89 : r_data = 29'b00000000000000000000000000000;
            8'h8A : r_data = 29'b00000000000000000000000000000;
            8'h8B : r_data = 29'b00000000000000000000000000000;
            8'h8C : r_data = 29'b00000000000000000000000000000;
            8'h8D : r_data = 29'b00000000000000000000000000000;
            8'h8E : r_data = 29'b00000000000000000000000000000;
            8'h8F : r_data = 29'b00000000000000000000000000000;
				
				//INC ACC
            8'h90 : r_data = 29'b11100011111110100001111000000;
            8'h91 : r_data = 29'b00000000000000000000000000000;
            8'h92 : r_data = 29'b00000000000000000000000000000;
            8'h93 : r_data = 29'b00000000000000000000000000000;
            8'h94 : r_data = 29'b00000000000000000000000000000;
            8'h95 : r_data = 29'b00000000000000000000000000000;
            8'h96 : r_data = 29'b00000000000000000000000000000;
            8'h97 : r_data = 29'b00000000000000000000000000000;
				
				//NEG ACC (CA2 ACC)         -- preguntar si lo vamos a poner 
            8'h98 : r_data = 29'b11110011111110000001111000000;  //este esta muy raro yo creo que no lo vamos a usar
            8'h99 : r_data = 29'b00000000000000000000000000000;
            8'h9A : r_data = 29'b00000000000000000000000000000;
            8'h9B : r_data = 29'b00000000000000000000000000000;
            8'h9C : r_data = 29'b00000000000000000000000000000;
            8'h9D : r_data = 29'b00000000000000000000000000000;
            8'h9E : r_data = 29'b00000000000000000000000000000;
            8'h9F : r_data = 29'b00000000000000000000000000000;
				
				//SLL ACC 
            8'hA0 : r_data = 29'b10001011111110100001111000000;
            8'hA1 : r_data = 29'b00000000000000000000000000000;
            8'hA2 : r_data = 29'b00000000000000000000000000000;
            8'hA3 : r_data = 29'b00000000000000000000000000000;
            8'hA4 : r_data = 29'b00000000000000000000000000000;
            8'hA5 : r_data = 29'b00000000000000000000000000000;
            8'hA6 : r_data = 29'b00000000000000000000000000000;
            8'hA7 : r_data = 29'b00000000000000000000000000000;
				
				//SLR ACC
            8'hA8 : r_data = 29'b10000111111110000001111000000;
            8'hA9 : r_data = 29'b00000000000000000000000000000;
            8'hAA : r_data = 29'b00000000000000000000000000000;
            8'hAB : r_data = 29'b00000000000000000000000000000;
            8'hAC : r_data = 29'b00000000000000000000000000000;
            8'hAD : r_data = 29'b00000000000000000000000000000;
            8'hAE : r_data = 29'b00000000000000000000000000000;
            8'hAF : r_data = 29'b00000000000000000000000000000;
				
				//CA2 ACC
            8'hB0 : r_data = 29'b11110011111110000001111000000;
            8'hB1 : r_data = 29'b00000000000000000000000000000;
            8'hB2 : r_data = 29'b00000000000000000000000000000;
            8'hB3 : r_data = 29'b00000000000000000000000000000;
            8'hB4 : r_data = 29'b00000000000000000000000000000;
            8'hB5 : r_data = 29'b00000000000000000000000000000;
            8'hB6 : r_data = 29'b00000000000000000000000000000;
            8'hB7 : r_data = 29'b00000000000000000000000000000;
				
				//SWAP ACC, A
            8'hB8 : r_data = 29'b10000001110110000000010000000;
            8'hB9 : r_data = 29'b00000011101110000000010000000;
            8'hBA : r_data = 29'b10000010111110000001111000000;
            8'hBB : r_data = 29'b00000000000000000000000000000;
            8'hBC : r_data = 29'b00000000000000000000000000000;
            8'hBD : r_data = 29'b00000000000000000000000000000;
            8'hBE : r_data = 29'b00000000000000000000000000000;
            8'hBF : r_data = 29'b00000000000000000000000000000;
				
				//MOV   DPTR, CTE

				
				8'hC0 : r_data = 29'b00000000000001000000010000000;
            8'hC1 : r_data = 29'b01100000000010000000010000000;
            8'hC2 : r_data = 29'b00000000000000110000010000000;
            8'hC3 : r_data = 29'b00000000001010010001111000000;
            8'hC4 : r_data = 29'b00000000000000000000000000000;
            8'hC5 : r_data = 29'b00000000000000000000000000000;
            8'hC6 : r_data = 29'b00000000000000000000000000000;
            8'hC7 : r_data = 29'b00000000000000000000000000000;
				
				//TODO ESTO DISPONIBLE PARA MAS INST...
            8'hC8 : r_data = 29'b00000000000000000000000000000;
            8'hC9 : r_data = 29'b00000000000000000000000000000;
            8'hCA : r_data = 29'b00000000000000000000000000000;
            8'hCB : r_data = 29'b00000000000000000000000000000;
            8'hCC : r_data = 29'b00000000000000000000000000000;
            8'hCD : r_data = 29'b00000000000000000000000000000;
            8'hCE : r_data = 29'b00000000000000000000000000000;
            8'hCF : r_data = 29'b00000000000000000000000000000;
				
				
            8'hD0 : r_data = 29'b00000000000000000000000000000;
            8'hD1 : r_data = 29'b00000000000000000000000000000;
            8'hD2 : r_data = 29'b00000000000000000000000000000;
            8'hD3 : r_data = 29'b00000000000000000000000000000;
            8'hD4 : r_data = 29'b00000000000000000000000000000;
            8'hD5 : r_data = 29'b00000000000000000000000000000;
            8'hD6 : r_data = 29'b00000000000000000000000000000;
            8'hD7 : r_data = 29'b00000000000000000000000000000;
            8'hD8 : r_data = 29'b00000000000000000000000000000;
            8'hD9 : r_data = 29'b00000000000000000000000000000;
            8'hDA : r_data = 29'b00000000000000000000000000000;
            8'hDB : r_data = 29'b00000000000000000000000000000;
            8'hDC : r_data = 29'b00000000000000000000000000000;
            8'hDD : r_data = 29'b00000000000000000000000000000;
            8'hDE : r_data = 29'b00000000000000000000000000000;
            8'hDF : r_data = 29'b00000000000000000000000000000;
            8'hE0 : r_data = 29'b00000000000000000000000000000;
            8'hE1 : r_data = 29'b00000000000000000000000000000;
            8'hE2 : r_data = 29'b00000000000000000000000000000;
            8'hE3 : r_data = 29'b00000000000000000000000000000;
            8'hE4 : r_data = 29'b00000000000000000000000000000;
            8'hE5 : r_data = 29'b00000000000000000000000000000;
            8'hE6 : r_data = 29'b00000000000000000000000000000;
            8'hE7 : r_data = 29'b00000000000000000000000000000;
            8'hE8 : r_data = 29'b00000000000000000000000000000;
            8'hE9 : r_data = 29'b00000000000000000000000000000;
            8'hEA : r_data = 29'b00000000000000000000000000000;
            8'hEB : r_data = 29'b00000000000000000000000000000;
            8'hEC : r_data = 29'b00000000000000000000000000000;
            8'hED : r_data = 29'b00000000000000000000000000000;
            8'hEE : r_data = 29'b00000000000000000000000000000;
            8'hEF : r_data = 29'b00000000000000000000000000000;
            8'hF0 : r_data = 29'b00000000000000000000000000000;
            8'hF1 : r_data = 29'b00000000000000000000000000000;
            8'hF2 : r_data = 29'b00000000000000000000000000000;
            8'hF3 : r_data = 29'b00000000000000000000000000000;
            8'hF4 : r_data = 29'b00000000000000000000000000000;
            8'hF5 : r_data = 29'b00000000000000000000000000000;
            8'hF6 : r_data = 29'b00000000000000000000000000000;
            8'hF7 : r_data = 29'b00000000000000000000000000000;
				
				//HALT
            8'hF8 : r_data = 29'b00000000000000000001111000000;
            8'hF9 : r_data = 29'b00000000000000000000000000000;
            8'hFA : r_data = 29'b00000000000000000000000000000;
            8'hFB : r_data = 29'b00000000000000000000000000000;
            8'hFC : r_data = 29'b00000000000000000000000000000;
            8'hFD : r_data = 29'b00000000000000000000000000000;
            8'hFE : r_data = 29'b00000000000000000000000000000;
            8'hFF : r_data = 29'b00000000000000000000000000000;
            default: r_data = 29'b00000000000000000000000000000;
        endcase

endmodule
